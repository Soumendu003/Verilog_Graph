module cf_ldpc_103(i1, i2, i3, o1);
  input [1:0] i1, i2, i3;
  output [1:0] o1;
  wire [1:0] i1, i2, i3;
  wire [1:0] o1;
  MX2X1 g35(.A (i3[1]), .B (i2[1]), .S0 (i1[1]), .Y (o1[1]));
  MX2X1 g36(.A (i3[0]), .B (i2[0]), .S0 (i1[0]), .Y (o1[0]));
endmodule

module cf_ldpc_102(i1, i2, i3, o1);
  input [2:0] i1, i2, i3;
  output [2:0] o1;
  wire [2:0] i1, i2, i3;
  wire [2:0] o1;
  cf_ldpc_103 s9(i1[1:0], i2[1:0], i3[1:0], o1[1:0]);
  MX2X1 g18(.A (i3[2]), .B (i2[2]), .S0 (i1[2]), .Y (o1[2]));
endmodule

module cf_ldpc_101(i1, i2, i3, o1);
  input [3:0] i1, i2, i3;
  output [3:0] o1;
  wire [3:0] i1, i2, i3;
  wire [3:0] o1;
  cf_ldpc_102 s9(i1[2:0], i2[2:0], i3[2:0], o1[2:0]);
  MX2X1 g18(.A (i3[3]), .B (i2[3]), .S0 (i1[3]), .Y (o1[3]));
endmodule

module cf_ldpc_100(i1, i2, i3, o1);
  input [4:0] i1, i2, i3;
  output [4:0] o1;
  wire [4:0] i1, i2, i3;
  wire [4:0] o1;
  cf_ldpc_101 s9(i1[3:0], i2[3:0], i3[3:0], o1[3:0]);
  MX2X1 g18(.A (i3[4]), .B (i2[4]), .S0 (i1[4]), .Y (o1[4]));
endmodule

module cf_ldpc_99(i1, i2, i3, o1);
  input [5:0] i1, i2, i3;
  output [5:0] o1;
  wire [5:0] i1, i2, i3;
  wire [5:0] o1;
  cf_ldpc_100 s9(i1[4:0], i2[4:0], i3[4:0], o1[4:0]);
  MX2X1 g18(.A (i3[5]), .B (i2[5]), .S0 (i1[5]), .Y (o1[5]));
endmodule

module cf_ldpc_98(i1, i2, i3, o1);
  input [6:0] i1, i2, i3;
  output [6:0] o1;
  wire [6:0] i1, i2, i3;
  wire [6:0] o1;
  cf_ldpc_99 s9(i1[5:0], i2[5:0], i3[5:0], o1[5:0]);
  MX2X1 g18(.A (i3[6]), .B (i2[6]), .S0 (i1[6]), .Y (o1[6]));
endmodule

module cf_ldpc_97(i1, i2, i3, o1);
  input [7:0] i1, i2, i3;
  output [7:0] o1;
  wire [7:0] i1, i2, i3;
  wire [7:0] o1;
  cf_ldpc_98 s9(i1[6:0], i2[6:0], i3[6:0], o1[6:0]);
  MX2X1 g18(.A (i3[7]), .B (i2[7]), .S0 (i1[7]), .Y (o1[7]));
endmodule

module cf_ldpc_96(i1, i2, i3, o1);
  input [8:0] i1, i2, i3;
  output [8:0] o1;
  wire [8:0] i1, i2, i3;
  wire [8:0] o1;
  cf_ldpc_97 s9(i1[7:0], i2[7:0], i3[7:0], o1[7:0]);
  MX2X1 g18(.A (i3[8]), .B (i2[8]), .S0 (i1[8]), .Y (o1[8]));
endmodule

module cf_ldpc_95(i1, i2, i3, o1);
  input [9:0] i1, i2, i3;
  output [9:0] o1;
  wire [9:0] i1, i2, i3;
  wire [9:0] o1;
  cf_ldpc_96 s9(i1[8:0], i2[8:0], i3[8:0], o1[8:0]);
  MX2X1 g18(.A (i3[9]), .B (i2[9]), .S0 (i1[9]), .Y (o1[9]));
endmodule

module cf_ldpc_94(i1, i2, i3, o1);
  input [10:0] i1, i2, i3;
  output [10:0] o1;
  wire [10:0] i1, i2, i3;
  wire [10:0] o1;
  cf_ldpc_95 s9(i1[9:0], i2[9:0], i3[9:0], o1[9:0]);
  MX2X1 g18(.A (i3[10]), .B (i2[10]), .S0 (i1[10]), .Y (o1[10]));
endmodule

module cf_ldpc_93(i1, i2, i3, o1);
  input [11:0] i1, i2, i3;
  output [11:0] o1;
  wire [11:0] i1, i2, i3;
  wire [11:0] o1;
  cf_ldpc_94 s9(i1[10:0], i2[10:0], i3[10:0], o1[10:0]);
  MX2X1 g18(.A (i3[11]), .B (i2[11]), .S0 (i1[11]), .Y (o1[11]));
endmodule

module cf_ldpc_92(i1, i2, i3, o1);
  input [12:0] i1, i2, i3;
  output [12:0] o1;
  wire [12:0] i1, i2, i3;
  wire [12:0] o1;
  cf_ldpc_93 s9(i1[11:0], i2[11:0], i3[11:0], o1[11:0]);
  MX2X1 g18(.A (i3[12]), .B (i2[12]), .S0 (i1[12]), .Y (o1[12]));
endmodule

module cf_ldpc_91(i1, i2, i3, o1);
  input [13:0] i1, i2, i3;
  output [13:0] o1;
  wire [13:0] i1, i2, i3;
  wire [13:0] o1;
  cf_ldpc_92 s9(i1[12:0], i2[12:0], i3[12:0], o1[12:0]);
  MX2X1 g18(.A (i3[13]), .B (i2[13]), .S0 (i1[13]), .Y (o1[13]));
endmodule

module cf_ldpc_90(i1, i2, i3, o1);
  input [14:0] i1, i2, i3;
  output [14:0] o1;
  wire [14:0] i1, i2, i3;
  wire [14:0] o1;
  cf_ldpc_91 s9(i1[13:0], i2[13:0], i3[13:0], o1[13:0]);
  MX2X1 g18(.A (i3[14]), .B (i2[14]), .S0 (i1[14]), .Y (o1[14]));
endmodule

module cf_ldpc_89(i1, i2, i3, o1);
  input [15:0] i1, i2, i3;
  output [15:0] o1;
  wire [15:0] i1, i2, i3;
  wire [15:0] o1;
  cf_ldpc_90 s9(i1[14:0], i2[14:0], i3[14:0], o1[14:0]);
  MX2X1 g18(.A (i3[15]), .B (i2[15]), .S0 (i1[15]), .Y (o1[15]));
endmodule

module cf_ldpc_88(i1, i2, i3, o1);
  input [16:0] i1, i2, i3;
  output [16:0] o1;
  wire [16:0] i1, i2, i3;
  wire [16:0] o1;
  cf_ldpc_89 s9(i1[15:0], i2[15:0], i3[15:0], o1[15:0]);
  MX2X1 g18(.A (i3[16]), .B (i2[16]), .S0 (i1[16]), .Y (o1[16]));
endmodule

module cf_ldpc_87(i1, i2, i3, o1);
  input [17:0] i1, i2, i3;
  output [17:0] o1;
  wire [17:0] i1, i2, i3;
  wire [17:0] o1;
  cf_ldpc_88 s9(i1[16:0], i2[16:0], i3[16:0], o1[16:0]);
  MX2X1 g18(.A (i3[17]), .B (i2[17]), .S0 (i1[17]), .Y (o1[17]));
endmodule

module cf_ldpc_86(i1, i2, i3, o1);
  input [18:0] i1, i2, i3;
  output [18:0] o1;
  wire [18:0] i1, i2, i3;
  wire [18:0] o1;
  cf_ldpc_87 s9(i1[17:0], i2[17:0], i3[17:0], o1[17:0]);
  MX2X1 g18(.A (i3[18]), .B (i2[18]), .S0 (i1[18]), .Y (o1[18]));
endmodule

module cf_ldpc_85(i1, i2, i3, o1);
  input [19:0] i1, i2, i3;
  output [19:0] o1;
  wire [19:0] i1, i2, i3;
  wire [19:0] o1;
  cf_ldpc_86 s9(i2[18:0], i3[18:0], i1[18:0], o1[18:0]);
  MX2X1 g17(.A (i1[19]), .B (i3[19]), .S0 (i2[19]), .Y (o1[19]));
endmodule

module cf_ldpc_84(i1, o1);
  input [19:0] i1;
  output o1;
  wire [19:0] i1;
  wire o1;
  wire n_0, n_1;
  OAI21X1 g19(.A0 (i1[5]), .A1 (n_0), .B0 (n_1), .Y (o1));
  NAND2XL g20(.A (i1[5]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_83(i1, o1);
  input [19:0] i1;
  output [1:0] o1;
  wire [19:0] i1;
  wire [1:0] o1;
  wire n_0, n_1;
  cf_ldpc_84 s10({4'b0000, i1[15], 4'b0000, i1[10], 4'b0000, i1[5],
       5'b00000}, o1[0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[1]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[8]), .B (i1[12]), .Y (n_0));
endmodule

module cf_ldpc_82(i1, o1);
  input [19:0] i1;
  output [2:0] o1;
  wire [19:0] i1;
  wire [2:0] o1;
  wire n_0, n_1;
  cf_ldpc_83 s10({4'b0000, i1[15], 2'b00, i1[12], 1'b0, i1[10], 1'b0,
       i1[8], 2'b00, i1[5:4], 4'b0000}, o1[1:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[2]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[2]), .B (i1[3]), .Y (n_0));
endmodule

module cf_ldpc_81(i1, o1);
  input [19:0] i1;
  output [3:0] o1;
  wire [19:0] i1;
  wire [3:0] o1;
  wire n_0, n_1;
  cf_ldpc_82 s10({4'b0000, i1[15], 2'b00, i1[12], 1'b0, i1[10], 1'b0,
       i1[8], 2'b00, i1[5:1], 1'b0}, o1[2:0]);
  OAI21X1 g19(.A0 (i1[7]), .A1 (n_0), .B0 (n_1), .Y (o1[3]));
  NAND2XL g20(.A (i1[7]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[12]), .B (i1[17]), .Y (n_0));
endmodule

module cf_ldpc_80(i1, o1);
  input [19:0] i1;
  output [4:0] o1;
  wire [19:0] i1;
  wire [4:0] o1;
  wire n_0, n_1;
  cf_ldpc_81 s10({2'b00, i1[17], 1'b0, i1[15], 2'b00, i1[12], 1'b0,
       i1[10], 1'b0, i1[8:7], 1'b0, i1[5:1], 1'b0}, o1[3:0]);
  OAI21X1 g19(.A0 (i1[5]), .A1 (n_0), .B0 (n_1), .Y (o1[4]));
  NAND2XL g20(.A (i1[5]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[16]), .B (i1[9]), .Y (n_0));
endmodule

module cf_ldpc_79(i1, o1);
  input [19:0] i1;
  output [5:0] o1;
  wire [19:0] i1;
  wire [5:0] o1;
  wire n_0, n_1;
  cf_ldpc_80 s10({2'b00, i1[17:15], 2'b00, i1[12], 1'b0, i1[10:7],
       1'b0, i1[5:1], 1'b0}, o1[4:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[5]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[2]), .B (i1[3]), .Y (n_0));
endmodule

module cf_ldpc_78(i1, o1);
  input [19:0] i1;
  output [6:0] o1;
  wire [19:0] i1;
  wire [6:0] o1;
  wire n_0, n_1;
  cf_ldpc_79 s10({2'b00, i1[17:15], 2'b00, i1[12], 1'b0, i1[10:7],
       1'b0, i1[5:0]}, o1[5:0]);
  OAI21X1 g19(.A0 (i1[8]), .A1 (n_0), .B0 (n_1), .Y (o1[6]));
  NAND2XL g20(.A (i1[8]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_77(i1, o1);
  input [19:0] i1;
  output [7:0] o1;
  wire [19:0] i1;
  wire [7:0] o1;
  wire n_0, n_1;
  cf_ldpc_78 s10({i1[19], 1'b0, i1[17:14], 1'b0, i1[12], 1'b0,
       i1[10:7], 1'b0, i1[5:0]}, o1[6:0]);
  OAI21X1 g19(.A0 (i1[6]), .A1 (n_0), .B0 (n_1), .Y (o1[7]));
  NAND2XL g20(.A (i1[6]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[13]), .B (i1[17]), .Y (n_0));
endmodule

module cf_ldpc_76(i1, o1);
  input [19:0] i1;
  output [8:0] o1;
  wire [19:0] i1;
  wire [8:0] o1;
  wire n_0, n_1;
  cf_ldpc_77 s10({i1[19], 1'b0, i1[17:12], 1'b0, i1[10:0]}, o1[7:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[8]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[1]), .B (i1[3]), .Y (n_0));
endmodule

module cf_ldpc_75(i1, o1);
  input [19:0] i1;
  output [9:0] o1;
  wire [19:0] i1;
  wire [9:0] o1;
  wire n_0, n_1;
  cf_ldpc_76 s10({i1[19], 1'b0, i1[17:12], 1'b0, i1[10:0]}, o1[8:0]);
  OAI21X1 g19(.A0 (i1[6]), .A1 (n_0), .B0 (n_1), .Y (o1[9]));
  NAND2XL g20(.A (i1[6]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[16]), .B (i1[11]), .Y (n_0));
endmodule

module cf_ldpc_74(i1, o1);
  input [19:0] i1;
  output [10:0] o1;
  wire [19:0] i1;
  wire [10:0] o1;
  wire n_0, n_1;
  cf_ldpc_75 s10({i1[19], 1'b0, i1[17:0]}, o1[9:0]);
  OAI21X1 g19(.A0 (i1[10]), .A1 (n_0), .B0 (n_1), .Y (o1[10]));
  NAND2XL g20(.A (i1[10]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[18]), .Y (n_0));
endmodule

module cf_ldpc_73(i1, o1);
  input [19:0] i1;
  output [11:0] o1;
  wire [19:0] i1;
  wire [11:0] o1;
  wire n_0, n_1;
  cf_ldpc_74 s10(i1, o1[10:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[11]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[1]), .B (i1[2]), .Y (n_0));
endmodule

module cf_ldpc_72(i1, o1);
  input [19:0] i1;
  output [12:0] o1;
  wire [19:0] i1;
  wire [12:0] o1;
  wire n_0, n_1;
  cf_ldpc_73 s10(i1, o1[11:0]);
  OAI21X1 g19(.A0 (i1[9]), .A1 (n_0), .B0 (n_1), .Y (o1[12]));
  NAND2XL g20(.A (i1[9]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[13]), .B (i1[18]), .Y (n_0));
endmodule

module cf_ldpc_71(i1, o1);
  input [19:0] i1;
  output [13:0] o1;
  wire [19:0] i1;
  wire [13:0] o1;
  wire n_0, n_1;
  cf_ldpc_72 s10(i1, o1[12:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[13]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[8]), .B (i1[12]), .Y (n_0));
endmodule

module cf_ldpc_70(i1, o1);
  input [19:0] i1;
  output [14:0] o1;
  wire [19:0] i1;
  wire [14:0] o1;
  wire n_0, n_1;
  cf_ldpc_71 s10(i1, o1[13:0]);
  OAI21X1 g19(.A0 (i1[5]), .A1 (n_0), .B0 (n_1), .Y (o1[14]));
  NAND2XL g20(.A (i1[5]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[6]), .B (i1[7]), .Y (n_0));
endmodule

module cf_ldpc_69(i1, o1);
  input [19:0] i1;
  output [15:0] o1;
  wire [19:0] i1;
  wire [15:0] o1;
  wire n_0, n_1;
  cf_ldpc_70 s10(i1, o1[14:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[15]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_68(i1, o1);
  input [19:0] i1;
  output [16:0] o1;
  wire [19:0] i1;
  wire [16:0] o1;
  wire n_0, n_1;
  cf_ldpc_69 s10(i1, o1[15:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[16]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[16]), .B (i1[9]), .Y (n_0));
endmodule

module cf_ldpc_67(i1, o1);
  input [19:0] i1;
  output [17:0] o1;
  wire [19:0] i1;
  wire [17:0] o1;
  wire n_0, n_1;
  cf_ldpc_68 s10(i1, o1[16:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[17]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[7]), .B (i1[6]), .Y (n_0));
endmodule

module cf_ldpc_66(i1, o1);
  input [19:0] i1;
  output [18:0] o1;
  wire [19:0] i1;
  wire [18:0] o1;
  wire n_0, n_1;
  cf_ldpc_67 s10(i1, o1[17:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[18]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[11]), .B (i1[16]), .Y (n_0));
endmodule

module cf_ldpc_65(i1, o1);
  input [19:0] i1;
  output [19:0] o1;
  wire [19:0] i1;
  wire [19:0] o1;
  wire n_0, n_1;
  cf_ldpc_66 s10(i1, o1[18:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[19]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[13]), .B (i1[17]), .Y (n_0));
endmodule

module cf_ldpc_64(i1, o1);
  input [19:0] i1;
  output [20:0] o1;
  wire [19:0] i1;
  wire [20:0] o1;
  wire n_0, n_1;
  cf_ldpc_65 s10(i1, o1[19:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[20]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[5]), .B (i1[7]), .Y (n_0));
endmodule

module cf_ldpc_63(i1, o1);
  input [19:0] i1;
  output [21:0] o1;
  wire [19:0] i1;
  wire [21:0] o1;
  wire n_0, n_1;
  cf_ldpc_64 s10(i1, o1[20:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[21]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[12]), .B (i1[17]), .Y (n_0));
endmodule

module cf_ldpc_62(i1, o1);
  input [19:0] i1;
  output [22:0] o1;
  wire [19:0] i1;
  wire [22:0] o1;
  wire n_0, n_1;
  cf_ldpc_63 s10(i1, o1[21:0]);
  OAI21X1 g19(.A0 (i1[11]), .A1 (n_0), .B0 (n_1), .Y (o1[22]));
  NAND2XL g20(.A (i1[11]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[15]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_61(i1, o1);
  input [19:0] i1;
  output [23:0] o1;
  wire [19:0] i1;
  wire [23:0] o1;
  wire n_0, n_1;
  cf_ldpc_62 s10(i1, o1[22:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[23]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[5]), .B (i1[6]), .Y (n_0));
endmodule

module cf_ldpc_60(i1, o1);
  input [19:0] i1;
  output [24:0] o1;
  wire [19:0] i1;
  wire [24:0] o1;
  wire n_0, n_1;
  cf_ldpc_61 s10(i1, o1[23:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[24]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_59(i1, o1);
  input [19:0] i1;
  output [25:0] o1;
  wire [19:0] i1;
  wire [25:0] o1;
  wire n_0, n_1;
  cf_ldpc_60 s10(i1, o1[24:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[25]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[4]), .B (i1[12]), .Y (n_0));
endmodule

module cf_ldpc_58(i1, o1);
  input [19:0] i1;
  output [26:0] o1;
  wire [19:0] i1;
  wire [26:0] o1;
  wire n_0, n_1;
  cf_ldpc_59 s10(i1, o1[25:0]);
  OAI21X1 g19(.A0 (i1[9]), .A1 (n_0), .B0 (n_1), .Y (o1[26]));
  NAND2XL g20(.A (i1[9]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[11]), .Y (n_0));
endmodule

module cf_ldpc_57(i1, o1);
  input [19:0] i1;
  output [27:0] o1;
  wire [19:0] i1;
  wire [27:0] o1;
  wire n_0, n_1;
  cf_ldpc_58 s10(i1, o1[26:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[27]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[18]), .B (i1[13]), .Y (n_0));
endmodule

module cf_ldpc_56(i1, o1);
  input [19:0] i1;
  output [28:0] o1;
  wire [19:0] i1;
  wire [28:0] o1;
  wire n_0, n_1;
  cf_ldpc_57 s10(i1, o1[27:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[28]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[16]), .B (i1[5]), .Y (n_0));
endmodule

module cf_ldpc_55(i1, o1);
  input [19:0] i1;
  output [29:0] o1;
  wire [19:0] i1;
  wire [29:0] o1;
  wire n_0, n_1;
  cf_ldpc_56 s10(i1, o1[28:0]);
  OAI21X1 g19(.A0 (i1[8]), .A1 (n_0), .B0 (n_1), .Y (o1[29]));
  NAND2XL g20(.A (i1[8]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[11]), .Y (n_0));
endmodule

module cf_ldpc_54(i1, o1);
  input [19:0] i1;
  output [30:0] o1;
  wire [19:0] i1;
  wire [30:0] o1;
  wire n_0, n_1;
  cf_ldpc_55 s10(i1, o1[29:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[30]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[15]), .B (i1[5]), .Y (n_0));
endmodule

module cf_ldpc_53(i1, o1);
  input [19:0] i1;
  output [31:0] o1;
  wire [19:0] i1;
  wire [31:0] o1;
  wire n_0, n_1;
  cf_ldpc_54 s10(i1, o1[30:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[31]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[18]), .Y (n_0));
endmodule

module cf_ldpc_52(i1, o1);
  input [19:0] i1;
  output [32:0] o1;
  wire [19:0] i1;
  wire [32:0] o1;
  wire n_0, n_1;
  cf_ldpc_53 s10(i1, o1[31:0]);
  OAI21X1 g19(.A0 (i1[8]), .A1 (n_0), .B0 (n_1), .Y (o1[32]));
  NAND2XL g20(.A (i1[8]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[9]), .B (i1[11]), .Y (n_0));
endmodule

module cf_ldpc_51(i1, o1);
  input [19:0] i1;
  output [33:0] o1;
  wire [19:0] i1;
  wire [33:0] o1;
  wire n_0, n_1;
  cf_ldpc_52 s10(i1, o1[32:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[33]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[16]), .B (i1[6]), .Y (n_0));
endmodule

module cf_ldpc_50(i1, o1);
  input [19:0] i1;
  output [34:0] o1;
  wire [19:0] i1;
  wire [34:0] o1;
  wire n_0, n_1;
  cf_ldpc_51 s10(i1, o1[33:0]);
  OAI21X1 g19(.A0 (i1[7]), .A1 (n_0), .B0 (n_1), .Y (o1[34]));
  NAND2XL g20(.A (i1[7]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[15]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_49(i1, o1);
  input [19:0] i1;
  output [35:0] o1;
  wire [19:0] i1;
  wire [35:0] o1;
  wire n_0, n_1;
  cf_ldpc_50 s10(i1, o1[34:0]);
  OAI21X1 g19(.A0 (i1[8]), .A1 (n_0), .B0 (n_1), .Y (o1[35]));
  NAND2XL g20(.A (i1[8]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[9]), .B (i1[10]), .Y (n_0));
endmodule

module cf_ldpc_48(i1, o1);
  input [19:0] i1;
  output [36:0] o1;
  wire [19:0] i1;
  wire [36:0] o1;
  wire n_0, n_1;
  cf_ldpc_49 s10(i1, o1[35:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[36]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[17]), .B (i1[7]), .Y (n_0));
endmodule

module cf_ldpc_47(i1, o1);
  input [19:0] i1;
  output [37:0] o1;
  wire [19:0] i1;
  wire [37:0] o1;
  wire n_0, n_1;
  cf_ldpc_48 s10(i1, o1[36:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[37]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[4]), .B (i1[8]), .Y (n_0));
endmodule

module cf_ldpc_46(i1, o1);
  input [19:0] i1;
  output [38:0] o1;
  wire [19:0] i1;
  wire [38:0] o1;
  wire n_0, n_1;
  cf_ldpc_47 s10(i1, o1[37:0]);
  OAI21X1 g19(.A0 (i1[13]), .A1 (n_0), .B0 (n_1), .Y (o1[38]));
  NAND2XL g20(.A (i1[13]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_45(i1, o1);
  input [19:0] i1;
  output [39:0] o1;
  wire [19:0] i1;
  wire [39:0] o1;
  wire n_0, n_1;
  cf_ldpc_46 s10(i1, o1[38:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[39]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[18]), .B (i1[9]), .Y (n_0));
endmodule

module cf_ldpc_44(i1, o1);
  input [19:0] i1;
  output [40:0] o1;
  wire [19:0] i1;
  wire [40:0] o1;
  wire n_0, n_1;
  cf_ldpc_45 s10(i1, o1[39:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[40]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[6]), .B (i1[17]), .Y (n_0));
endmodule

module cf_ldpc_43(i1, o1);
  input [19:0] i1;
  output [41:0] o1;
  wire [19:0] i1;
  wire [41:0] o1;
  wire n_0, n_1;
  cf_ldpc_44 s10(i1, o1[40:0]);
  OAI21X1 g19(.A0 (i1[12]), .A1 (n_0), .B0 (n_1), .Y (o1[41]));
  NAND2XL g20(.A (i1[12]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[14]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_42(i1, o1);
  input [19:0] i1;
  output [42:0] o1;
  wire [19:0] i1;
  wire [42:0] o1;
  wire n_0, n_1;
  cf_ldpc_43 s10(i1, o1[41:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[42]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[19]), .B (i1[8]), .Y (n_0));
endmodule

module cf_ldpc_41(i1, o1);
  input [19:0] i1;
  output [43:0] o1;
  wire [19:0] i1;
  wire [43:0] o1;
  wire n_0, n_1;
  cf_ldpc_42 s10(i1, o1[42:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[43]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[18]), .Y (n_0));
endmodule

module cf_ldpc_40(i1, o1);
  input [19:0] i1;
  output [44:0] o1;
  wire [19:0] i1;
  wire [44:0] o1;
  wire n_0, n_1;
  cf_ldpc_41 s10(i1, o1[43:0]);
  OAI21X1 g19(.A0 (i1[12]), .A1 (n_0), .B0 (n_1), .Y (o1[44]));
  NAND2XL g20(.A (i1[12]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[13]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_39(i1, o1);
  input [19:0] i1;
  output [45:0] o1;
  wire [19:0] i1;
  wire [45:0] o1;
  wire n_0, n_1;
  cf_ldpc_40 s10(i1, o1[44:0]);
  OAI21X1 g19(.A0 (i1[0]), .A1 (n_0), .B0 (n_1), .Y (o1[45]));
  NAND2XL g20(.A (i1[0]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[5]), .B (i1[10]), .Y (n_0));
endmodule

module cf_ldpc_38(i1, o1);
  input [19:0] i1;
  output [46:0] o1;
  wire [19:0] i1;
  wire [46:0] o1;
  wire n_0, n_1;
  cf_ldpc_39 s10(i1, o1[45:0]);
  OAI21X1 g19(.A0 (i1[7]), .A1 (n_0), .B0 (n_1), .Y (o1[46]));
  NAND2XL g20(.A (i1[7]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[11]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_37(i1, o1);
  input [19:0] i1;
  output [47:0] o1;
  wire [19:0] i1;
  wire [47:0] o1;
  wire n_0, n_1;
  cf_ldpc_38 s10(i1, o1[46:0]);
  OAI21X1 g19(.A0 (i1[12]), .A1 (n_0), .B0 (n_1), .Y (o1[47]));
  NAND2XL g20(.A (i1[12]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[13]), .B (i1[14]), .Y (n_0));
endmodule

module cf_ldpc_36(i1, o1);
  input [19:0] i1;
  output [48:0] o1;
  wire [19:0] i1;
  wire [48:0] o1;
  wire n_0, n_1;
  cf_ldpc_37 s10(i1, o1[47:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[48]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[6]), .B (i1[11]), .Y (n_0));
endmodule

module cf_ldpc_35(i1, o1);
  input [19:0] i1;
  output [49:0] o1;
  wire [19:0] i1;
  wire [49:0] o1;
  wire n_0, n_1;
  cf_ldpc_36 s10(i1, o1[48:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[49]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[5]), .B (i1[9]), .Y (n_0));
endmodule

module cf_ldpc_34(i1, o1);
  input [19:0] i1;
  output [50:0] o1;
  wire [19:0] i1;
  wire [50:0] o1;
  wire n_0, n_1;
  cf_ldpc_35 s10(i1, o1[49:0]);
  OAI21X1 g19(.A0 (i1[17]), .A1 (n_0), .B0 (n_1), .Y (o1[50]));
  NAND2XL g20(.A (i1[17]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[18]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_33(i1, o1);
  input [19:0] i1;
  output [51:0] o1;
  wire [19:0] i1;
  wire [51:0] o1;
  wire n_0, n_1;
  cf_ldpc_34 s10(i1, o1[50:0]);
  OAI21X1 g19(.A0 (i1[1]), .A1 (n_0), .B0 (n_1), .Y (o1[51]));
  NAND2XL g20(.A (i1[1]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[12]), .B (i1[7]), .Y (n_0));
endmodule

module cf_ldpc_32(i1, o1);
  input [19:0] i1;
  output [52:0] o1;
  wire [19:0] i1;
  wire [52:0] o1;
  wire n_0, n_1;
  cf_ldpc_33 s10(i1, o1[51:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[52]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[6]), .B (i1[13]), .Y (n_0));
endmodule

module cf_ldpc_31(i1, o1);
  input [19:0] i1;
  output [53:0] o1;
  wire [19:0] i1;
  wire [53:0] o1;
  wire n_0, n_1;
  cf_ldpc_32 s10(i1, o1[52:0]);
  OAI21X1 g19(.A0 (i1[16]), .A1 (n_0), .B0 (n_1), .Y (o1[53]));
  NAND2XL g20(.A (i1[16]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[18]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_30(i1, o1);
  input [19:0] i1;
  output [54:0] o1;
  wire [19:0] i1;
  wire [54:0] o1;
  wire n_0, n_1;
  cf_ldpc_31 s10(i1, o1[53:0]);
  OAI21X1 g27(.A0 (i1[4]), .A1 (n_0), .B0 (n_1), .Y (o1[54]));
  NAND2XL g28(.A (i1[4]), .B (n_0), .Y (n_1));
  XNOR2X1 g29(.A (i1[9]), .B (i1[13]), .Y (n_0));
endmodule

module cf_ldpc_29(i1, o1);
  input [19:0] i1;
  output [55:0] o1;
  wire [19:0] i1;
  wire [55:0] o1;
  wire n_0, n_1;
  cf_ldpc_30 s10(i1, o1[54:0]);
  OAI21X1 g19(.A0 (i1[3]), .A1 (n_0), .B0 (n_1), .Y (o1[55]));
  NAND2XL g20(.A (i1[3]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[10]), .B (i1[14]), .Y (n_0));
endmodule

module cf_ldpc_28(i1, o1);
  input [19:0] i1;
  output [56:0] o1;
  wire [19:0] i1;
  wire [56:0] o1;
  wire n_0, n_1;
  cf_ldpc_29 s10(i1, o1[55:0]);
  OAI21X1 g19(.A0 (i1[16]), .A1 (n_0), .B0 (n_1), .Y (o1[56]));
  NAND2XL g20(.A (i1[16]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[17]), .B (i1[19]), .Y (n_0));
endmodule

module cf_ldpc_27(i1, o1);
  input [19:0] i1;
  output [57:0] o1;
  wire [19:0] i1;
  wire [57:0] o1;
  wire n_0, n_1;
  cf_ldpc_28 s10(i1, o1[56:0]);
  OAI21X1 g19(.A0 (i1[2]), .A1 (n_0), .B0 (n_1), .Y (o1[57]));
  NAND2XL g20(.A (i1[2]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[8]), .B (i1[14]), .Y (n_0));
endmodule

module cf_ldpc_26(i1, o1);
  input [19:0] i1;
  output [58:0] o1;
  wire [19:0] i1;
  wire [58:0] o1;
  wire n_0, n_1;
  cf_ldpc_27 s10(i1, o1[57:0]);
  OAI21X1 g19(.A0 (i1[7]), .A1 (n_0), .B0 (n_1), .Y (o1[58]));
  NAND2XL g20(.A (i1[7]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[11]), .B (i1[15]), .Y (n_0));
endmodule

module cf_ldpc_25(i1, o1);
  input [19:0] i1;
  output [59:0] o1;
  wire [19:0] i1;
  wire [59:0] o1;
  wire n_0, n_1;
  cf_ldpc_26 s10(i1, o1[58:0]);
  OAI21X1 g19(.A0 (i1[16]), .A1 (n_0), .B0 (n_1), .Y (o1[59]));
  NAND2XL g20(.A (i1[16]), .B (n_0), .Y (n_1));
  XNOR2X1 g21(.A (i1[17]), .B (i1[18]), .Y (n_0));
endmodule

module cf_ldpc_21(i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12,
     i13, i14, i15, o1);
  input i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14,
       i15;
  output o1;
  wire i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15;
  wire o1;
  wire n_0, n_1, n_2, n_3;
  NAND4XL g93(.A (n_3), .B (n_2), .C (n_1), .D (n_0), .Y (o1));
  NOR3X1 g94(.A (i12), .B (i4), .C (i15), .Y (n_3));
  NOR4X1 g95(.A (i10), .B (i9), .C (i8), .D (i11), .Y (n_2));
  NOR4X1 g96(.A (i2), .B (i6), .C (i3), .D (i7), .Y (n_1));
  NOR4X1 g97(.A (i14), .B (i13), .C (i1), .D (i5), .Y (n_0));
endmodule

module cf_ldpc_20_14(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_11(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_0), .A1 (n_1), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_0), .B (n_1), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[0]), .B (i1[1]), .Y (n_0));
endmodule

module cf_ldpc_20_8(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_5(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  XNOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XOR2X1 g33(.A (i1[0]), .B (i1[1]), .Y (n_0));
endmodule

module cf_ldpc_20(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_1(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_2(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_19(i1, o1);
  input [19:0] i1;
  output [2:0] o1;
  wire [19:0] i1;
  wire [2:0] o1;
  cf_ldpc_20 s6({i1[15], i1[10], i1[5], i1[0]}, o1[0]);
  cf_ldpc_20_1 s7({i1[16], i1[11], i1[6], i1[3]}, o1[1]);
  cf_ldpc_20_2 s8({i1[17], i1[12], i1[7], i1[1]}, o1[2]);
endmodule

module cf_ldpc_20_3(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_0), .A1 (n_1), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_0), .B (n_1), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[0]), .B (i1[1]), .Y (n_0));
endmodule

module cf_ldpc_20_4(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_18(i1, o1);
  input [19:0] i1;
  output [5:0] o1;
  wire [19:0] i1;
  wire [5:0] o1;
  cf_ldpc_20_5 s10({i1[12], i1[8], i1[4], i1[0]}, o1[5]);
  cf_ldpc_19 s7({2'b00, i1[17:15], 2'b00, i1[12:10], 2'b00, i1[7:5],
       1'b0, i1[3], 1'b0, i1[1:0]}, o1[2:0]);
  cf_ldpc_20_3 s8({i1[18], i1[13], i1[9], i1[4]}, o1[3]);
  cf_ldpc_20_4 s9({i1[19], i1[14], i1[8], i1[2]}, o1[4]);
endmodule

module cf_ldpc_20_6(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_7(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_17(i1, o1);
  input [19:0] i1;
  output [8:0] o1;
  wire [19:0] i1;
  wire [8:0] o1;
  cf_ldpc_20_8 s10({i1[18], i1[14], i1[10], i1[3]}, o1[8]);
  cf_ldpc_18 s7(i1, o1[5:0]);
  cf_ldpc_20_6 s8({i1[16], i1[9], i1[5], i1[1]}, o1[6]);
  cf_ldpc_20_7 s9({i1[17], i1[13], i1[6], i1[2]}, o1[7]);
endmodule

module cf_ldpc_20_9(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_10(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_16(i1, o1);
  input [19:0] i1;
  output [11:0] o1;
  wire [19:0] i1;
  wire [11:0] o1;
  cf_ldpc_20_11 s10(i1[7:4], o1[11]);
  cf_ldpc_17 s7(i1, o1[8:0]);
  cf_ldpc_20_9 s8({i1[19], i1[15], i1[11], i1[7]}, o1[9]);
  cf_ldpc_20_10 s9(i1[3:0], o1[10]);
endmodule

module cf_ldpc_20_12(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_20_13(i1, o1);
  input [3:0] i1;
  output o1;
  wire [3:0] i1;
  wire o1;
  wire n_0, n_1, n_2;
  OAI21X1 g30(.A0 (n_1), .A1 (n_0), .B0 (n_2), .Y (o1));
  NAND2XL g31(.A (n_1), .B (n_0), .Y (n_2));
  CLKXOR2X1 g32(.A (i1[2]), .B (i1[3]), .Y (n_1));
  XNOR2X1 g33(.A (i1[1]), .B (i1[0]), .Y (n_0));
endmodule

module cf_ldpc_15(i1, o1);
  input [19:0] i1;
  output [14:0] o1;
  wire [19:0] i1;
  wire [14:0] o1;
  cf_ldpc_20_14 s10(i1[19:16], o1[14]);
  cf_ldpc_16 s7(i1, o1[11:0]);
  cf_ldpc_20_12 s8(i1[11:8], o1[12]);
  cf_ldpc_20_13 s9(i1[15:12], o1[13]);
endmodule

module cf_ldpc_14(i1, o1);
  input [19:0] i1;
  output o1;
  wire [19:0] i1;
  wire o1;
  wire [14:0] s8_1;
  wire s7_1;
  cf_ldpc_21 s7(s8_1[14], s8_1[13], s8_1[12], s8_1[11], s8_1[10],
       s8_1[9], s8_1[8], s8_1[7], s8_1[6], s8_1[5], s8_1[4], s8_1[3],
       s8_1[2], s8_1[1], s8_1[0], s7_1);
  cf_ldpc_15 s8(i1, s8_1);
  INVXL g2(.A (s7_1), .Y (o1));
endmodule

module cf_ldpc_13_18(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_18(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_18 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_16(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_16(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_16 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_14(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_14(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_14 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_12(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_12(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_12 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_10(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_10(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_10 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_8(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_8(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_8 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_6(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_6(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_6 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_4(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[0]), .B (i1[1]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_4(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_4 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_2(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_2(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_2 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13 s9(i1, s9_1);
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_13_1(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_1(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_1 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_11(i1, o1, o2);
  input [5:0] i1;
  output [1:0] o1, o2;
  wire [5:0] i1;
  wire [1:0] o1, o2;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  cf_ldpc_12 s7(i1[2:0], o1[0]);
  cf_ldpc_12_1 s8(i1[5:3], o1[1]);
endmodule

module cf_ldpc_13_3(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_3(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_3 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_10(i1, o1, o2);
  input [11:0] i1;
  output [3:0] o1, o2;
  wire [11:0] i1;
  wire [3:0] o1, o2;
  wire UNCONNECTED, UNCONNECTED0;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  cf_ldpc_12_2 s11(i1[8:6], o1[2]);
  cf_ldpc_11 s12(i1[5:0], o1[1:0], {UNCONNECTED0, UNCONNECTED});
  cf_ldpc_12_3 s13(i1[11:9], o1[3]);
endmodule

module cf_ldpc_13_5(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_5(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_5 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_9(i1, o1, o2);
  input [17:0] i1;
  output [5:0] o1, o2;
  wire [17:0] i1;
  wire [5:0] o1, o2;
  wire UNCONNECTED1, UNCONNECTED2, UNCONNECTED3, UNCONNECTED4;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  cf_ldpc_12_4 s11(i1[14:12], o1[4]);
  cf_ldpc_10 s12(i1[11:0], o1[3:0], {UNCONNECTED4, UNCONNECTED3,
       UNCONNECTED2, UNCONNECTED1});
  cf_ldpc_12_5 s13(i1[17:15], o1[5]);
endmodule

module cf_ldpc_13_7(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_7(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_7 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_8(i1, o1, o2);
  input [23:0] i1;
  output [7:0] o1, o2;
  wire [23:0] i1;
  wire [7:0] o1, o2;
  wire UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8,
       UNCONNECTED9, UNCONNECTED10;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  cf_ldpc_12_6 s11(i1[20:18], o1[6]);
  cf_ldpc_9 s12(i1[17:0], o1[5:0], {UNCONNECTED10, UNCONNECTED9,
       UNCONNECTED8, UNCONNECTED7, UNCONNECTED6, UNCONNECTED5});
  cf_ldpc_12_7 s13(i1[23:21], o1[7]);
endmodule

module cf_ldpc_13_9(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_9(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_9 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_7(i1, o1, o2);
  input [29:0] i1;
  output [9:0] o1, o2;
  wire [29:0] i1;
  wire [9:0] o1, o2;
  wire UNCONNECTED11, UNCONNECTED12, UNCONNECTED13, UNCONNECTED14,
       UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  cf_ldpc_12_8 s11(i1[26:24], o1[8]);
  cf_ldpc_8 s12(i1[23:0], o1[7:0], {UNCONNECTED18, UNCONNECTED17,
       UNCONNECTED16, UNCONNECTED15, UNCONNECTED14, UNCONNECTED13,
       UNCONNECTED12, UNCONNECTED11});
  cf_ldpc_12_9 s13(i1[29:27], o1[9]);
endmodule

module cf_ldpc_13_11(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_11(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_11 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_6(i1, o1, o2);
  input [35:0] i1;
  output [11:0] o1, o2;
  wire [35:0] i1;
  wire [11:0] o1, o2;
  wire UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22,
       UNCONNECTED23, UNCONNECTED24, UNCONNECTED25, UNCONNECTED26;
  wire UNCONNECTED27, UNCONNECTED28;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  assign o2[10] = 1'b0;
  assign o2[11] = 1'b0;
  cf_ldpc_12_10 s11(i1[32:30], o1[10]);
  cf_ldpc_7 s12(i1[29:0], o1[9:0], {UNCONNECTED28, UNCONNECTED27,
       UNCONNECTED26, UNCONNECTED25, UNCONNECTED24, UNCONNECTED23,
       UNCONNECTED22, UNCONNECTED21, UNCONNECTED20, UNCONNECTED19});
  cf_ldpc_12_11 s13(i1[35:33], o1[11]);
endmodule

module cf_ldpc_13_13(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_13(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_13 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_5(i1, o1, o2);
  input [41:0] i1;
  output [13:0] o1, o2;
  wire [41:0] i1;
  wire [13:0] o1, o2;
  wire UNCONNECTED29, UNCONNECTED30, UNCONNECTED31, UNCONNECTED32,
       UNCONNECTED33, UNCONNECTED34, UNCONNECTED35, UNCONNECTED36;
  wire UNCONNECTED37, UNCONNECTED38, UNCONNECTED39, UNCONNECTED40;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  assign o2[10] = 1'b0;
  assign o2[11] = 1'b0;
  assign o2[12] = 1'b0;
  assign o2[13] = 1'b0;
  cf_ldpc_12_12 s11(i1[38:36], o1[12]);
  cf_ldpc_6 s12(i1[35:0], o1[11:0], {UNCONNECTED40, UNCONNECTED39,
       UNCONNECTED38, UNCONNECTED37, UNCONNECTED36, UNCONNECTED35,
       UNCONNECTED34, UNCONNECTED33, UNCONNECTED32, UNCONNECTED31,
       UNCONNECTED30, UNCONNECTED29});
  cf_ldpc_12_13 s13(i1[41:39], o1[13]);
endmodule

module cf_ldpc_13_15(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_15(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_15 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_4(i1, o1, o2);
  input [47:0] i1;
  output [15:0] o1, o2;
  wire [47:0] i1;
  wire [15:0] o1, o2;
  wire UNCONNECTED41, UNCONNECTED42, UNCONNECTED43, UNCONNECTED44,
       UNCONNECTED45, UNCONNECTED46, UNCONNECTED47, UNCONNECTED48;
  wire UNCONNECTED49, UNCONNECTED50, UNCONNECTED51, UNCONNECTED52,
       UNCONNECTED53, UNCONNECTED54;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  assign o2[10] = 1'b0;
  assign o2[11] = 1'b0;
  assign o2[12] = 1'b0;
  assign o2[13] = 1'b0;
  assign o2[14] = 1'b0;
  assign o2[15] = 1'b0;
  cf_ldpc_12_14 s11(i1[44:42], o1[14]);
  cf_ldpc_5 s12(i1[41:0], o1[13:0], {UNCONNECTED54, UNCONNECTED53,
       UNCONNECTED52, UNCONNECTED51, UNCONNECTED50, UNCONNECTED49,
       UNCONNECTED48, UNCONNECTED47, UNCONNECTED46, UNCONNECTED45,
       UNCONNECTED44, UNCONNECTED43, UNCONNECTED42, UNCONNECTED41});
  cf_ldpc_12_15 s13(i1[47:45], o1[15]);
endmodule

module cf_ldpc_13_17(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_17(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_17 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_3(i1, o1, o2);
  input [53:0] i1;
  output [17:0] o1, o2;
  wire [53:0] i1;
  wire [17:0] o1, o2;
  wire UNCONNECTED55, UNCONNECTED56, UNCONNECTED57, UNCONNECTED58,
       UNCONNECTED59, UNCONNECTED60, UNCONNECTED61, UNCONNECTED62;
  wire UNCONNECTED63, UNCONNECTED64, UNCONNECTED65, UNCONNECTED66,
       UNCONNECTED67, UNCONNECTED68, UNCONNECTED69, UNCONNECTED70;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  assign o2[10] = 1'b0;
  assign o2[11] = 1'b0;
  assign o2[12] = 1'b0;
  assign o2[13] = 1'b0;
  assign o2[14] = 1'b0;
  assign o2[15] = 1'b0;
  assign o2[16] = 1'b0;
  assign o2[17] = 1'b0;
  cf_ldpc_12_16 s11(i1[50:48], o1[16]);
  cf_ldpc_4 s12(i1[47:0], o1[15:0], {UNCONNECTED70, UNCONNECTED69,
       UNCONNECTED68, UNCONNECTED67, UNCONNECTED66, UNCONNECTED65,
       UNCONNECTED64, UNCONNECTED63, UNCONNECTED62, UNCONNECTED61,
       UNCONNECTED60, UNCONNECTED59, UNCONNECTED58, UNCONNECTED57,
       UNCONNECTED56, UNCONNECTED55});
  cf_ldpc_12_17 s13(i1[53:51], o1[17]);
endmodule

module cf_ldpc_13_19(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  NOR3X1 g19(.A (i1[1]), .B (i1[0]), .C (i1[2]), .Y (o1));
endmodule

module cf_ldpc_12_19(i1, o1);
  input [2:0] i1;
  output o1;
  wire [2:0] i1;
  wire o1;
  wire n_0, s9_1;
  cf_ldpc_13_19 s9(.i1 (i1), .o1 (s9_1));
  CLKINVX1 g25(.A (n_0), .Y (o1));
  AOI31X1 g26(.A0 (i1[1]), .A1 (i1[0]), .A2 (i1[2]), .B0 (s9_1), .Y
       (n_0));
endmodule

module cf_ldpc_2(i1, o1, o2);
  input [59:0] i1;
  output [19:0] o1, o2;
  wire [59:0] i1;
  wire [19:0] o1, o2;
  wire UNCONNECTED71, UNCONNECTED72, UNCONNECTED73, UNCONNECTED74,
       UNCONNECTED75, UNCONNECTED76, UNCONNECTED77, UNCONNECTED78;
  wire UNCONNECTED79, UNCONNECTED80, UNCONNECTED81, UNCONNECTED82,
       UNCONNECTED83, UNCONNECTED84, UNCONNECTED85, UNCONNECTED86;
  wire UNCONNECTED87, UNCONNECTED88;
  assign o2[0] = 1'b0;
  assign o2[1] = 1'b0;
  assign o2[2] = 1'b0;
  assign o2[3] = 1'b0;
  assign o2[4] = 1'b0;
  assign o2[5] = 1'b0;
  assign o2[6] = 1'b0;
  assign o2[7] = 1'b0;
  assign o2[8] = 1'b0;
  assign o2[9] = 1'b0;
  assign o2[10] = 1'b0;
  assign o2[11] = 1'b0;
  assign o2[12] = 1'b0;
  assign o2[13] = 1'b0;
  assign o2[14] = 1'b0;
  assign o2[15] = 1'b0;
  assign o2[16] = 1'b0;
  assign o2[17] = 1'b0;
  assign o2[18] = 1'b0;
  assign o2[19] = 1'b0;
  cf_ldpc_12_18 s11(i1[56:54], o1[18]);
  cf_ldpc_3 s12(i1[53:0], o1[17:0], {UNCONNECTED88, UNCONNECTED87,
       UNCONNECTED86, UNCONNECTED85, UNCONNECTED84, UNCONNECTED83,
       UNCONNECTED82, UNCONNECTED81, UNCONNECTED80, UNCONNECTED79,
       UNCONNECTED78, UNCONNECTED77, UNCONNECTED76, UNCONNECTED75,
       UNCONNECTED74, UNCONNECTED73, UNCONNECTED72, UNCONNECTED71});
  cf_ldpc_12_19 s13(i1[59:57], o1[19]);
endmodule

module cf_ldpc_1(clock_c, i1, i2, o1, o2);
  input clock_c, i1;
  input [19:0] i2;
  output o1;
  output [19:0] o2;
  wire clock_c, i1;
  wire [19:0] i2;
  wire o1;
  wire [19:0] o2;
  wire [19:0] n3;
  wire [19:0] s9_1;
  wire [59:0] s7_1;
  wire [19:0] s6_1;
  wire UNCONNECTED89, UNCONNECTED90, UNCONNECTED91, UNCONNECTED92,
       UNCONNECTED93, UNCONNECTED94, UNCONNECTED95, UNCONNECTED96;
  wire UNCONNECTED97, UNCONNECTED98, UNCONNECTED99, UNCONNECTED100,
       UNCONNECTED101, UNCONNECTED102, UNCONNECTED103, UNCONNECTED104;
  wire UNCONNECTED105, UNCONNECTED106, UNCONNECTED107, UNCONNECTED108;
  cf_ldpc_85 s6(n3, s9_1, {s7_1[59], s7_1[56], s7_1[53], s7_1[50],
       s7_1[47], s7_1[44], s7_1[41], s7_1[38], s7_1[35], s7_1[32],
       s7_1[29], s7_1[26], s7_1[23], s7_1[20], s7_1[17], s7_1[14],
       s7_1[11], s7_1[8], s7_1[5], s7_1[2]}, s6_1);
  cf_ldpc_25 s7(o2, s7_1);
  cf_ldpc_14 s8(o2, o1);
  cf_ldpc_2 s9(s7_1, s9_1, {UNCONNECTED108, UNCONNECTED107,
       UNCONNECTED106, UNCONNECTED105, UNCONNECTED104, UNCONNECTED103,
       UNCONNECTED102, UNCONNECTED101, UNCONNECTED100, UNCONNECTED99,
       UNCONNECTED98, UNCONNECTED97, UNCONNECTED96, UNCONNECTED95,
       UNCONNECTED94, UNCONNECTED93, UNCONNECTED92, UNCONNECTED91,
       UNCONNECTED90, UNCONNECTED89});
  SDFFQX1 \n5_reg[4] (.CK (clock_c), .D (s6_1[4]), .SI (i2[4]), .SE
       (i1), .Q (o2[4]));
  SDFFQX1 \n3_reg[0] (.CK (clock_c), .D (n3[0]), .SI (i2[0]), .SE (i1),
       .Q (n3[0]));
  SDFFQX1 \n3_reg[10] (.CK (clock_c), .D (n3[10]), .SI (i2[10]), .SE
       (i1), .Q (n3[10]));
  SDFFQX1 \n3_reg[1] (.CK (clock_c), .D (n3[1]), .SI (i2[1]), .SE (i1),
       .Q (n3[1]));
  SDFFQX1 \n3_reg[2] (.CK (clock_c), .D (n3[2]), .SI (i2[2]), .SE (i1),
       .Q (n3[2]));
  SDFFQX1 \n3_reg[3] (.CK (clock_c), .D (n3[3]), .SI (i2[3]), .SE (i1),
       .Q (n3[3]));
  SDFFQX1 \n3_reg[4] (.CK (clock_c), .D (n3[4]), .SI (i2[4]), .SE (i1),
       .Q (n3[4]));
  SDFFQX1 \n3_reg[5] (.CK (clock_c), .D (n3[5]), .SI (i2[5]), .SE (i1),
       .Q (n3[5]));
  SDFFQX1 \n3_reg[6] (.CK (clock_c), .D (n3[6]), .SI (i2[6]), .SE (i1),
       .Q (n3[6]));
  SDFFQX1 \n3_reg[7] (.CK (clock_c), .D (n3[7]), .SI (i2[7]), .SE (i1),
       .Q (n3[7]));
  SDFFQX1 \n3_reg[8] (.CK (clock_c), .D (n3[8]), .SI (i2[8]), .SE (i1),
       .Q (n3[8]));
  SDFFQX1 \n3_reg[11] (.CK (clock_c), .D (n3[11]), .SI (i2[11]), .SE
       (i1), .Q (n3[11]));
  SDFFQX1 \n3_reg[9] (.CK (clock_c), .D (n3[9]), .SI (i2[9]), .SE (i1),
       .Q (n3[9]));
  SDFFQX1 \n5_reg[0] (.CK (clock_c), .D (s6_1[0]), .SI (i2[0]), .SE
       (i1), .Q (o2[0]));
  SDFFQX1 \n5_reg[10] (.CK (clock_c), .D (s6_1[10]), .SI (i2[10]), .SE
       (i1), .Q (o2[10]));
  SDFFQX1 \n5_reg[11] (.CK (clock_c), .D (s6_1[11]), .SI (i2[11]), .SE
       (i1), .Q (o2[11]));
  SDFFQX1 \n5_reg[12] (.CK (clock_c), .D (s6_1[12]), .SI (i2[12]), .SE
       (i1), .Q (o2[12]));
  SDFFQX1 \n5_reg[13] (.CK (clock_c), .D (s6_1[13]), .SI (i2[13]), .SE
       (i1), .Q (o2[13]));
  SDFFQX1 \n5_reg[14] (.CK (clock_c), .D (s6_1[14]), .SI (i2[14]), .SE
       (i1), .Q (o2[14]));
  SDFFQX1 \n5_reg[15] (.CK (clock_c), .D (s6_1[15]), .SI (i2[15]), .SE
       (i1), .Q (o2[15]));
  SDFFQX1 \n3_reg[12] (.CK (clock_c), .D (n3[12]), .SI (i2[12]), .SE
       (i1), .Q (n3[12]));
  SDFFQX1 \n3_reg[13] (.CK (clock_c), .D (n3[13]), .SI (i2[13]), .SE
       (i1), .Q (n3[13]));
  SDFFQX1 \n5_reg[16] (.CK (clock_c), .D (s6_1[16]), .SI (i2[16]), .SE
       (i1), .Q (o2[16]));
  SDFFQX1 \n5_reg[17] (.CK (clock_c), .D (s6_1[17]), .SI (i2[17]), .SE
       (i1), .Q (o2[17]));
  SDFFQX1 \n5_reg[18] (.CK (clock_c), .D (s6_1[18]), .SI (i2[18]), .SE
       (i1), .Q (o2[18]));
  SDFFQX1 \n5_reg[19] (.CK (clock_c), .D (s6_1[19]), .SI (i2[19]), .SE
       (i1), .Q (o2[19]));
  SDFFQX1 \n3_reg[14] (.CK (clock_c), .D (n3[14]), .SI (i2[14]), .SE
       (i1), .Q (n3[14]));
  SDFFQX1 \n5_reg[1] (.CK (clock_c), .D (s6_1[1]), .SI (i2[1]), .SE
       (i1), .Q (o2[1]));
  SDFFQX1 \n5_reg[2] (.CK (clock_c), .D (s6_1[2]), .SI (i2[2]), .SE
       (i1), .Q (o2[2]));
  SDFFQX1 \n3_reg[15] (.CK (clock_c), .D (n3[15]), .SI (i2[15]), .SE
       (i1), .Q (n3[15]));
  SDFFQX1 \n5_reg[3] (.CK (clock_c), .D (s6_1[3]), .SI (i2[3]), .SE
       (i1), .Q (o2[3]));
  SDFFQX1 \n5_reg[5] (.CK (clock_c), .D (s6_1[5]), .SI (i2[5]), .SE
       (i1), .Q (o2[5]));
  SDFFQX1 \n3_reg[16] (.CK (clock_c), .D (n3[16]), .SI (i2[16]), .SE
       (i1), .Q (n3[16]));
  SDFFQX1 \n3_reg[17] (.CK (clock_c), .D (n3[17]), .SI (i2[17]), .SE
       (i1), .Q (n3[17]));
  SDFFQX1 \n5_reg[6] (.CK (clock_c), .D (s6_1[6]), .SI (i2[6]), .SE
       (i1), .Q (o2[6]));
  SDFFQX1 \n5_reg[7] (.CK (clock_c), .D (s6_1[7]), .SI (i2[7]), .SE
       (i1), .Q (o2[7]));
  SDFFQX1 \n5_reg[8] (.CK (clock_c), .D (s6_1[8]), .SI (i2[8]), .SE
       (i1), .Q (o2[8]));
  SDFFQX1 \n5_reg[9] (.CK (clock_c), .D (s6_1[9]), .SI (i2[9]), .SE
       (i1), .Q (o2[9]));
  SDFFQX1 \n3_reg[18] (.CK (clock_c), .D (n3[18]), .SI (i2[18]), .SE
       (i1), .Q (n3[18]));
  SDFFQX1 \n3_reg[19] (.CK (clock_c), .D (n3[19]), .SI (i2[19]), .SE
       (i1), .Q (n3[19]));
endmodule

module cf_ldpc(clock_c, start_i, message_i, valid_o, message_o);
  input clock_c, start_i;
  input [19:0] message_i;
  output valid_o;
  output [19:0] message_o;
  wire clock_c, start_i;
  wire [19:0] message_i;
  wire valid_o;
  wire [19:0] message_o;
  cf_ldpc_1 s1(clock_c, start_i, message_i, valid_o, message_o);
endmodule

